library IEEE;
use IEEE.STD_LOGIC_1164.all;

package Utility is
	 TYPE myArray is ARRAY (natural range <>) OF STD_LOGIC_VECTOR(15 DOWNTO 0);
	 TYPE myArray2D is array (natural range <>, natural range <>) of std_logic_vector(15 downto 0);
end Utility;

package body Utility is
end Utility;
